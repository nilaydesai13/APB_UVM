`include "uvm_macros.svh"

package apb_pkg;
	import uvm_pkg::*;
	`include "apb_master_trans.sv"
	`include "apb_seq.sv"
	`include "apb_sequencer.sv"
	`include "apb_master_driver.sv"
	`include "apb_monitor.sv"
	`include "apb_agent.sv"
	`include "apb_scoreboard.sv"
	`include "apb_env.sv"
	`include "apb_test.sv"
endpackage